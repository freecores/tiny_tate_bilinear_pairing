/*
    Copyright 2012 Homer Hsing
    
    This file is part of Tiny Tate Bilinear Pairing Core.

    Tiny Tate Bilinear Pairing Core is free software: you can redistribute it and/or modify
    it under the terms of the GNU Lesser General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    Tiny Tate Bilinear Pairing Core is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU Lesser General Public License for more details.

    You should have received a copy of the GNU Lesser General Public License
    along with Tiny Tate Bilinear Pairing Core.  If not, see http://www.gnu.org/licenses/lgpl.txt
*/

module rom (clk, addr, out);
   input clk;
   input [8:0] addr;
   output reg [28:0] out;
   
   always @(posedge clk)
      case (addr)
         0: out <= 29'h1860042;
         1: out <= 29'h30d0041;
         2: out <= 29'h38f0041;
         3: out <= 29'h60046;
         4: out <= 29'hb01b180;
         5: out <= 29'hb810041;
         6: out <= 29'hb8bb197;
         7: out <= 29'hc0bb187;
         8: out <= 29'hcb1b187;
         9: out <= 29'h7ae8059;
         10: out <= 29'h79e8045;
         11: out <= 29'hbb1b185;
         12: out <= 29'hc2fb180;
         13: out <= 29'hb0fb196;
         14: out <= 29'h8b00056;
         15: out <= 29'h8a20051;
         16: out <= 29'h90a0045;
         17: out <= 29'h98fb180;
         18: out <= 29'h9ae8053;
         19: out <= 29'ha020041;
         20: out <= 29'ha8e0047;
         21: out <= 29'h1f0041;
         22: out <= 29'hb230041;
         23: out <= 29'hba50041;
         24: out <= 29'hc270041;
         25: out <= 29'hca90041;
         26: out <= 29'hd2b0041;
         27: out <= 29'h7800057;
         28: out <= 29'h79e0059;
         29: out <= 29'h8ac0058;
         30: out <= 29'h8a2005a;
         31: out <= 29'h8a20051;
         32: out <= 29'h92e8059;
         33: out <= 29'h9b48058;
         34: out <= 29'ha320041;
         35: out <= 29'hab4005a;
         36: out <= 29'h30d0081;
         37: out <= 29'h30c8042;
         38: out <= 29'h38f0081;
         39: out <= 29'h38e0047;
         40: out <= 29'h60046;
         41: out <= 29'hb000040;
         42: out <= 29'hb8bb187;
         43: out <= 29'h2db180;
         44: out <= 29'hc000056;
         45: out <= 29'hc808056;
         46: out <= 29'hd1e0054;
         47: out <= 29'hdb40052;
         48: out <= 29'he348052;
         49: out <= 29'he9e8054;
         50: out <= 29'hf3a8053;
         51: out <= 29'heba0053;
         52: out <= 29'hfa20055;
         53: out <= 29'h103e0053;
         54: out <= 29'h10be8053;
         55: out <= 29'h112e0056;
         56: out <= 29'hb2e8056;
         57: out <= 29'h11a28055;
         58: out <= 29'h12460052;
         59: out <= 29'h11c68052;
         60: out <= 29'h12b00057;
         61: out <= 29'h13360060;
         62: out <= 29'h13800062;
         63: out <= 29'h143c0064;
         64: out <= 29'h14b20057;
         65: out <= 29'h15380061;
         66: out <= 29'h15800056;
         67: out <= 29'h163a0063;
         68: out <= 29'hc31b19b;
         69: out <= 29'hdcbb1a6;
         70: out <= 29'h102fb1a0;
         71: out <= 29'hf01b19e;
         72: out <= 29'h12cfb1a8;
         73: out <= 29'h1145b1a4;
         74: out <= 29'hcb3b19c;
         75: out <= 29'he53b1aa;
         76: out <= 29'hbafb1a1;
         77: out <= 29'h1b19d;
         78: out <= 29'hed7b1ac;
         79: out <= 29'hb2db1a3;
         80: out <= 29'h10b00065;
         81: out <= 29'h11c0005d;
         82: out <= 29'h12408057;
         83: out <= 29'h13328058;
         84: out <= 29'hbae0060;
         85: out <= 29'hbc48057;
         86: out <= 29'hbae0056;
         87: out <= 29'hc320058;
         88: out <= 29'hc30805e;
         89: out <= 29'hc308040;
         90: out <= 29'hcc68061;
         91: out <= 29'hcb2805e;
         92: out <= 29'hb320056;
         93: out <= 29'hcc20063;
         94: out <= 29'hcb2805b;
         95: out <= 29'hcb20062;
         96: out <= 29'h320040;
         97: out <= 29'hcc80066;
         98: out <= 29'hf488066;
         99: out <= 29'hf3c005c;
         100: out <= 29'hf3c805b;
         101: out <= 29'h102e0058;
         102: out <= 29'hbae8058;
         103: out <= 29'hbae005c;
         104: out <= 29'hbae005b;
         105: out <= 29'hbae8065;
         106: out <= 29'hbae805d;
         107: out <= 29'h7ac8052;
         108: out <= 29'h8808053;
         109: out <= 29'h328052;
         110: out <= 29'h8054;
         111: out <= 29'hb3c8053;
         112: out <= 29'hb2c8055;
         113: out <= 29'ha40805a;
         114: out <= 29'haae805f;
         115: out <= 29'h9008041;
         116: out <= 29'h9ac8041;
         117: out <= 29'h49f0041;
         118: out <= 29'h1e0052;
         119: out <= 29'h54;
         120: out <= 29'hb1fb18f;
         121: out <= 29'hb9fb192;
         122: out <= 29'hc25b194;
         123: out <= 29'hca9b194;
         124: out <= 29'h1b180;
         125: out <= 29'hbae0058;
         126: out <= 29'hc2c8058;
         127: out <= 29'hcb28057;
         128: out <= 29'h57;
         129: out <= 29'h8056;
         130: out <= 29'hb220053;
         131: out <= 29'hb2c0055;
         132: out <= 29'hba3b191;
         133: out <= 29'hd23b193;
         134: out <= 29'hda7b195;
         135: out <= 29'he2bb195;
         136: out <= 29'hb2db196;
         137: out <= 29'hd34005b;
         138: out <= 29'hdae805b;
         139: out <= 29'he38805a;
         140: out <= 29'hb2c005a;
         141: out <= 29'hb2c8057;
         142: out <= 29'hb9e0052;
         143: out <= 29'hd1e0054;
         144: out <= 29'hea40054;
         145: out <= 29'hf220053;
         146: out <= 29'hfa20055;
         147: out <= 29'h10260055;
         148: out <= 29'h109fb191;
         149: out <= 29'h1125b193;
         150: out <= 29'h11a9b195;
         151: out <= 29'hbafb19e;
         152: out <= 29'hd35b19f;
         153: out <= 29'hebbb1a0;
         154: out <= 29'hf428062;
         155: out <= 29'hfbc8063;
         156: out <= 29'hfbe005d;
         157: out <= 29'hbae805e;
         158: out <= 29'hbae005d;
         159: out <= 29'hd34805e;
         160: out <= 29'heb0805b;
         161: out <= 29'hf32805c;
         162: out <= 29'h10008056;
         163: out <= 29'hc30005b;
         164: out <= 29'hcb2005c;
         165: out <= 29'h56;
         166: out <= 29'hb300059;
         167: out <= 29'hdb08040;
         168: out <= 29'he328058;
         169: out <= 29'h1080805c;
         170: out <= 29'h1131b198;
         171: out <= 29'h11b3b199;
         172: out <= 29'h1201b180;
         173: out <= 29'hcb1b199;
         174: out <= 29'hc31b180;
         175: out <= 29'h1b196;
         176: out <= 29'hb45b19b;
         177: out <= 29'hdc7b19c;
         178: out <= 29'he49b1a1;
         179: out <= 29'hb2c005b;
         180: out <= 29'hb2c005c;
         181: out <= 29'hdac0041;
         182: out <= 29'he370041;
         183: out <= 29'he37b19c;
         184: out <= 29'h10b90041;
         185: out <= 29'hdb7b1a1;
         186: out <= 29'h10b70081;
         187: out <= 29'he39b1a1;
         188: out <= 29'h10b900c1;
         189: out <= 29'hdb7b1a1;
         190: out <= 29'h10b70201;
         191: out <= 29'hdb7b1a1;
         192: out <= 29'h10b70141;
         193: out <= 29'he39b1a1;
         194: out <= 29'he390401;
         195: out <= 29'hdb7b19c;
         196: out <= 29'he370941;
         197: out <= 29'hdb7b19c;
         198: out <= 29'he371281;
         199: out <= 29'hdb7b19c;
         200: out <= 29'he372501;
         201: out <= 29'hdb7b19c;
         202: out <= 29'he374a01;
         203: out <= 29'hdb7b19c;
         204: out <= 29'hdb70041;
         205: out <= 29'hb37b196;
         206: out <= 29'hb37b196;
         207: out <= 29'hdc68064;
         208: out <= 29'he44805b;
         209: out <= 29'h388040;
         210: out <= 29'hcc88059;
         211: out <= 29'hc368058;
         212: out <= 29'h2db180;
         213: out <= 29'hcadb199;
         214: out <= 29'hb2db198;
         215: out <= 29'hc3a005e;
         216: out <= 29'hdba0060;
         217: out <= 29'he3c0060;
         218: out <= 29'h10800059;
         219: out <= 29'h11000056;
         220: out <= 29'h11b20056;
         221: out <= 29'hebbb180;
         222: out <= 29'hf3db199;
         223: out <= 29'h1041b196;
         224: out <= 29'hc31b1a1;
         225: out <= 29'hdb7b1a2;
         226: out <= 29'he39b1a3;
         227: out <= 29'heba805e;
         228: out <= 29'hf3a8060;
         229: out <= 29'hf3c005c;
         230: out <= 29'hc30805d;
         231: out <= 29'hc30005c;
         232: out <= 29'hdb6805d;
         233: out <= 29'he3e0057;
         234: out <= 29'hebe005a;
         235: out <= 29'h102e005a;
         236: out <= 29'h10800059;
         237: out <= 29'h11000056;
         238: out <= 29'h11b20056;
         239: out <= 29'h3fb180;
         240: out <= 29'hbafb199;
         241: out <= 29'hb35b196;
         242: out <= 29'hcb9b1a1;
         243: out <= 29'hd3bb1a2;
         244: out <= 29'he41b1a3;
         245: out <= 29'h8057;
         246: out <= 29'hb008056;
         247: out <= 29'hb2c005c;
         248: out <= 29'hbb28040;
         249: out <= 29'hbae005c;
         250: out <= 29'h348040;
         251: out <= 29'hcbc0056;
         252: out <= 29'hd300057;
         253: out <= 29'he368040;
         254: out <= 29'hebdb19b;
         255: out <= 29'hfadb180;
         256: out <= 29'hdb1b19b;
         257: out <= 29'h2fb180;
         258: out <= 29'h1033b19c;
         259: out <= 29'hb2db198;
         260: out <= 29'hbbdb197;
         261: out <= 29'hc33b19a;
         262: out <= 29'hcb5b19c;
         263: out <= 29'hd2c0057;
         264: out <= 29'hc348058;
         265: out <= 29'hd360040;
         266: out <= 29'hd34005a;
         267: out <= 29'h805b;
         268: out <= 29'hdbe805d;
         269: out <= 29'hdb60060;
         270: out <= 29'he04005d;
         271: out <= 29'he38005f;
         272: out <= 29'he38805a;
         273: out <= 29'hb2e8056;
         274: out <= 29'hb360056;
         275: out <= 29'hbb00041;
         276: out <= 29'heb20040;
         277: out <= 29'hdba005b;
         278: out <= 29'hc30005a;
         279: out <= 29'hc300058;
         280: out <= 29'h320040;
         281: out <= 29'h40;
         282: out <= 29'hcb90041;
         283: out <= 29'hd2d0041;
         284: out <= 29'heaf0041;
         285: out <= 29'hf370041;
         286: out <= 29'hfb10041;
         287: out <= 29'h10010041;
         288: out <= 29'hcb2005d;
         289: out <= 29'hcb2005f;
         290: out <= 29'hd34005a;
         291: out <= 29'hd34805e;
         292: out <= 29'hd348060;
         293: out <= 29'heba805f;
         294: out <= 29'hf40805e;
         295: out <= 29'h10400060;
         296: out <= 29'hcb30041;
         297: out <= 29'hd350041;
         298: out <= 29'hebb0041;
         299: out <= 29'hf3d0041;
         300: out <= 29'hfbf0041;
         301: out <= 29'h10410041;
         302: out <= 29'hcb2005d;
         303: out <= 29'hcb2005f;
         304: out <= 29'hd34005a;
         305: out <= 29'hd34805e;
         306: out <= 29'hd348060;
         307: out <= 29'heba805f;
         308: out <= 29'hf40805e;
         309: out <= 29'h10400060;
         310: out <= 29'h10b80056;
         311: out <= 29'h112e005b;
         312: out <= 29'h11b08040;
         313: out <= 29'h1239b198;
         314: out <= 29'h12adb180;
         315: out <= 29'hc2fb198;
         316: out <= 29'h37b180;
         317: out <= 29'h1343b1a3;
         318: out <= 29'hb2db197;
         319: out <= 29'hbb9b19b;
         320: out <= 29'hdc3b1a2;
         321: out <= 29'he45b1a3;
         322: out <= 29'h10ac0057;
         323: out <= 29'hdc2805b;
         324: out <= 29'h10b00040;
         325: out <= 29'h10c20061;
         326: out <= 29'h8058;
         327: out <= 29'hc4a8064;
         328: out <= 29'hc300066;
         329: out <= 29'h11040064;
         330: out <= 29'h11440065;
         331: out <= 29'h11448061;
         332: out <= 29'hb2e8056;
         333: out <= 29'hb300056;
         334: out <= 29'hbb60041;
         335: out <= 29'h11b80040;
         336: out <= 29'hc460058;
         337: out <= 29'hdb60061;
         338: out <= 29'hdb6005b;
         339: out <= 29'h380040;
         340: out <= 29'h40;
         341: out <= 29'he32005f;
         342: out <= 29'h10b8005d;
         343: out <= 29'he38805d;
         344: out <= 29'h11c4005b;
         345: out <= 29'h12460057;
         346: out <= 29'h11c68057;
         347: out <= 29'hcb2805f;
         348: out <= 29'h12b2805e;
         349: out <= 29'hcb2005e;
         350: out <= 29'h1144805b;
         351: out <= 29'h13448058;
         352: out <= 29'h11440058;
         353: out <= 29'h13b40060;
         354: out <= 29'h144e005e;
         355: out <= 29'hf4e805e;
         356: out <= 29'h13ac0040;
         357: out <= 29'h14ce0058;
         358: out <= 29'hc4e8058;
         359: out <= 29'hd348060;
         360: out <= 29'h13b4005d;
         361: out <= 29'hd34805d;
         362: out <= 29'hb2c8040;
         363: out <= 29'heac0057;
         364: out <= 29'hb2c8057;
         365: out <= 29'hbc20068;
         366: out <= 29'h15480069;
         367: out <= 29'h15ca0067;
         368: out <= 29'h164c005d;
         369: out <= 29'h16b8005e;
         370: out <= 29'h17460058;
         371: out <= 29'h17b2005a;
         372: out <= 29'h18440056;
         373: out <= 29'h18be0060;
         374: out <= 29'h19360040;
         375: out <= 29'h10c3b1a4;
         376: out <= 29'hbafb1aa;
         377: out <= 29'h1251b1a9;
         378: out <= 29'h12cbb1a6;
         379: out <= 29'h1357b1ac;
         380: out <= 29'hecfb19d;
         381: out <= 29'he39b1a3;
         382: out <= 29'h11dbb1ae;
         383: out <= 29'hc3db198;
         384: out <= 29'hcb3b1a2;
         385: out <= 29'hf5fb1b0;
         386: out <= 29'hb35b196;
         387: out <= 29'hd3fb19b;
         388: out <= 29'hde3b1b2;
         389: out <= 29'h41b180;
         390: out <= 29'hfc20066;
         391: out <= 29'hfbe005a;
         392: out <= 29'h1048005e;
         393: out <= 29'h10400040;
         394: out <= 29'hd38005a;
         395: out <= 29'h300040;
         396: out <= 29'h40;
         397: out <= 29'hc46005b;
         398: out <= 29'he000064;
         399: out <= 29'h11348061;
         400: out <= 29'h8064;
         401: out <= 29'h5d;
         402: out <= 29'h56;
         403: out <= 29'hd340061;
         404: out <= 29'hd348065;
         405: out <= 29'hd348059;
         406: out <= 29'h4c0805f;
         407: out <= 29'h4928065;
         408: out <= 29'h4920056;
         409: out <= 29'h53e0060;
         410: out <= 29'h5148057;
         411: out <= 29'h514005d;
         412: out <= 29'h5140059;
         413: out <= 29'h514805b;
         414: out <= 29'h5b80062;
         415: out <= 29'h6388062;
         416: out <= 29'h6180058;
         417: out <= 29'h6188057;
         418: out <= 29'h680005a;
         419: out <= 29'h700805a;
         420: out <= 29'h71c0058;
         421: out <= 29'h71c0057;
         422: out <= 29'h71c8066;
         423: out <= 29'h71c805e;
         default: out <= 0;
      endcase
endmodule
